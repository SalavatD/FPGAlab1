`timescale 1ns / 1ps

// ������ ������������ ������ main:
module main_tb(

    );
    
    ///////////////////////////////////////////// ���������� //////////////////////////////////////
    
    reg  [9:0] sw;      // 10-�� ��������� ����
    wire [9:0] led;     // ����� LED �����������
    wire [6:0] hex;     // ����� �� 7-�� ���������� ���������
    wire [7:0] hex_on;  // ����� ��� ���������� ��������� ������������
    
    // ����������� ���������� ������ main:
    main DUT (
    .sw     (sw),
    .led    (led),
    .hex    (hex),
    .hex_on (hex_on)
    );
    
    ///////////////////////////////////////////// ����������� ��� /////////////////////////////////
    
    initial begin
        // ������ SW[9:8] = 00
        // �� DC-DEC ��������� ����� DC1
        sw = 10'b0;
        #5 sw[3:0] = 4'b1;
        #5 sw[3:0] = 4'b11;
        #5 sw[3:0] = 4'b111;
        #5 sw[3:0] = 4'b1111;
        
        // ������ SW[9:8] = 01
        // �� DC-DEC ��������� ����� DC2
        #5 sw[3:0] = 8'h0;
        sw[7:4] = 4'b0;
        sw[9:8] = 2'b1;
        #5 sw[7:4] = 4'b0010;
        #5 sw[7:4] = 4'b1101;
        #5 sw[7:4] = 4'b1111;
        
        // ������ SW[9:8] = 10
        // �� DC-DEC ��������� ����� �������
        #5 sw[7:0] = 8'h0;
        sw[9:8] = 2'b10;
        #5 sw[3:0] = 4'b0101;
        #5 sw[3:0] = 4'b1010;
        #5 sw[3:0] = 4'b1111;
        
        // ������ SW[9:8] = 11
        // �� DC-DEC ��������� SW[3:0]
        #5 sw[7:0] = 8'h0;
        sw[9:8] = 2'b11;
        #5 sw[3:0] = 4'h1;
        #5 sw[3:0] = 4'h2;
        #5 sw[3:0] = 4'h3;
        #5 sw[3:0] = 4'h4;
        #5 sw[3:0] = 4'h5;
        #5 sw[3:0] = 4'h6;
        #5 sw[3:0] = 4'h7;
        #5 sw[3:0] = 4'h8;
        #5 sw[3:0] = 4'h9;
        #5 sw[3:0] = 4'hA;
        #5 sw[3:0] = 4'hB;
        #5 sw[3:0] = 4'hC;
        #5 sw[3:0] = 4'hD;
        #5 sw[3:0] = 4'hE;
        #5 sw[3:0] = 4'hF;
        #5 $stop;
    end
    
endmodule
